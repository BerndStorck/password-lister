UILANG="Svenska"
LABEL_PASSWORD_FILE="Lösenordsfil"

ERROR="FEL"
ERR_MISSING_CONFIGURATION_FILE="Ingen konfigurationsfil hittades!"
THE_FILE="Filen"
NOT_FOUND="hittades inte"

WARNING="VARNING"
DISALLOWED_OPTION="Otillåtet alternativ"
